BY FABRIZIO CARUSO LEVEL COMPLETED GAME COMPETED CROSS BOMBER NEW HISCORE DESTROY ALL PRESS FIRE GAME OVER BUILDINGS LEVEL BONUS joy���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ����L ` 0�cL:��� � mc�� 0��  .穠 �� ��e�f g�c��	� �� ��g�h�d�d��L7��� � mc�� �� 0�d .�0 �� �� 0��  .��� p� ���	�H�@e	�h 0�g�hmd���i��	� � �   ��� � mc�� �� 0�d .�0 �� �� 0��  .��� p� �����	�H�@e	�h 0�g�hmd���i��	� � à  ���dLU��c g�c��	��L�L�� 0�i�i�� �L�� F�
 _�j� �j �� F�
 � �� �� �q �� ��8�iH�� �h 0��  .穠 �� ��l�m� �j�0 ��  ��n�o�k�k��L�¢ �� �q �� ��8�iH�� �h �� 0�k .�0 �� �� 0��  .��� p� ���	�H�@e	�h 0�n�omk���i��	� � �   �� �� �q �� ��8�iH�� �h �� 0�k .�0 �� �� 0��  .��� p� �����	�H�@e	�h 0�n�omk���i��	� � à  ���kL���iLT�L� � � �@��	� �@ �� L�� � � JJJJ���	� �L�� � )���	� � �L�� 0� g��	��L%Ġ i��	� � ��q�r�p�p��LĠ� � 
�� 0�p .�0 �� �� 0��  .��� p� ���	�H�@e	�h 0�q�rmp���i��	� � �   ��� � 
�� 0�p .�0 �� �� 0��  .��� p� �����	�H�@e	�h 0�q�rmp���i��	� � à  ���pLC� g��	� L�Ĝs�t�t� ��s��L�Ġ� � 
�� 0�s�t 0�0 �� �� 0��  .��� p� ���	���@e	�	� ���� 
�� 0�s�t 0�0 �� �� 0��  .��� p� �����	���@e	�	� ��s�L+��tL+� g��	��L�`�u�u��`�v�v��L�Ŝw�x�x� ��w��L�Ţ �u
�� 0�w�x 0�0 �� �� 0�v .��� p� ���	���@e	�	� ���u
�� 0�w�x 0�0 �� �� 0�v .��� p� �����	���@e	�	� ��w�L��xL��vL���uL�ĩ  N) �� N) ��` 0� .� i� �� ��J ��  � i� �L�� ��U� 札�������������� X� �ĩ �1�� �ũ � �� �ũ �J�� �ũ	 �k�� �ũ �V�� ��L�ᜣ������������ �ĩ � �u�� �� � � � �� N� �� �Ĝ�����L�Ǣ �! �䍵��������L�Ǣ ��
�� 0筴 .�0 �� ���	��e��e	�	�H�@e	�h 0筵��m����i��	� � �   �� ��
�� 0筴 .�0 �� ���	��eH�e	�h���	�H�@e	�h 0筵��m����i��	� � à  ���L���L�Ɯ����� � ��
��iy��i�	� �����٩������LEɢ ��
��iy��i�� 0筦 .� � �� 0� n�) ��  �� n�)
����������� �� 0� ��
��iy��i�� Z� ��L?ɭ��	���� � �䍸����� ����L9ɭ�
�� 0筷 .�0 �� �� 0�8�H� � �h 0��� p� ���	�H�@e	�h 0筸��m����i��	� � �   �� ��
�� 0筷 .�0 �� �� 0�8�H� � �h 0��� p� �����	�H�@e	�h 0筸��m����i��	� � à  �� �LS��L��L�ǩ��:�� �  � 筧�� N�� �& �䍻����� ����L� .�0 ���	�H�@e	�h 0筻��m����i��	� � �   �筺 .�0 �����	�H�@e	�h 0筻��m����i��	� � à  �� �Lxɭ' �䍾����� ����L�� .�0 �� ���	�H�@e	�h 0签��m����i��	� � �   �筽 .�0 �� �����	�H�@e	�h 0签��m����i��	� � à  �� �Lʭ( �������� ����LQ� .�0 �� ���	�H�@e	�h 0����m����i��	� � �   ��� .�0 �� �����	�H�@e	�h 0����m����i��	� � à  �� ��L�ʭ) �����������L�˭� .�0 �� ���	�H�@e	�h 0����m����i��	� � �   ��� .�0 �� �����	�H�@e	�h 0����m����i��	� � à  ����L`˩ �  � � �� N�� �# �����������L�̭� .�0 �� ���	�H�@e	�h 0����m����i��	� � �   ��� .�0 �� �����	�H�@e	�h 0����m����i��	� � à  ����L̩	 �  � � �� N�� �  � 筭�� N�L�ݭ��Ljέ���Ljέ���LjΜ������ �����L�͢ �� �� �� 0���� 0�0 �� �� 0筢 .��� p� ���	���@e	�	� ���� �� �� 0���� 0�0 �� �� 0筢 .��� p� �����	���@e	�	� ����L���L͜������ �����Le΢ ��
�� 0���� 0�0 �� �� 0筢 .��� p� ���	���@e	�	� ����
�� 0���� 0�0 �� �� 0筢 .��� p� �����	���@e	�	� ����L����L���� � �������� ����LQϭ� �� �� 0�� .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0����m����i��	� � �   �� �� �� �� 0�� .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0����m����i��	� � à  �� ��L{έ �������� ����L4Э�
�� 0�� .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0����m����i��	� � �   �� ��
�� 0�� .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0����m����i��	� � à  �� ��Lbϭ �������� ����Lѭ��� �� 0�� .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0����m����i��	� � �   �� ���� �� 0�� .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0����m����i��	� � à  �� ��LEМ������� 0��� 0� �� � �� �� ��
�������ӭ��L�ҭ��LҜ������ �����LҢ ��
�� 0���� 0�0 �� �� 0筥 .��� p� ���	���@e	�	� ����
�� 0���� 0�0 �� �� 0筥 .��� p� �����	���@e	�	� ����Lf���Lfќ�����L`ש  N) �L`����������� ��
��iy��i�	���L`ע ��
��iy��i�	� ����
m�����ί�'�8�H� � �h �� 0筦 .� �� �䍩��� �  � 筧�� N�L`ע � �������� ����L�ӭ�
�� 0�� .�0 �� �� 0筥 .��� p� ���	�H�@e	�h 0����m����i��	� � �   �� ��
�� 0�� .�0 �� �� 0筥 .��� p� �����	�H�@e	�h 0����m����i��	� � à  �� ��L�ҭ  �����������L�Ԣ ��
�� 0�� .�0 �� �� 0� ���� 0��� p� ���	�H�@e	�h 0����m����i��	� � �   �� ��
�� 0�� .�0 �� �� 0� ���� 0��� p� �����	�H�@e	�h 0����m����i��	� � à  ����L������� �L`׭ �����������L�բ ��
�� 0�� .�0 �� �� 0筥 .��� p� ���	�H�@e	�h 0����m����i��	� � �   �� ��
�� 0�� .�0 �� �� 0筥 .��� p� �����	�H�@e	�h 0����m����i��	� � à  ����L�Ԝ�����	 �  � � �� N�������� �����L]֢ ��
�� 0���� 0�0 �� �� 0� �� �� 0��� p� ���	���@e	�	� ����
�� 0���� 0�0 �� �� 0� �� �� 0��� p� �����	���@e	�	� ����L����L�բ �* �������� ����LB׭�
�� 0�� .�0 �� �� 0筥 .��� p� ���	�H�@e	�h 0����m����i��	� � �   �� ��
�� 0�� .�0 �� �� 0筥 .��� p� �����	�H�@e	�h 0����m����i��	� � à  �� ��Lp֜����������c�
�������������� �����Lآ �� �� �� 0���� 0�0 �� �� 0筢 .��� p� ���	���@e	�	� ���� �� �� 0���� 0�0 �� �� 0筢 .��� p� �����	���@e	�	� ����Lf���Lfע � �������� ����L�ح�
�� 0�� .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0����m����i��	� � �   �� ��
�� 0�� .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0����m����i��	� � à  �� ��L%ح �������� ����L�٭��� �� 0�� .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0����m����i��	� � �   �� ���� �� 0�� .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0����m����i��	� � à  �� ��Lٜ������� 0��� 0� �� � �� �� ��
�������ӭ��L�ۢ � �������� ����L ۭ�
�� 0�� .�0 �� �� 0筥 .��� p� ���	�H�@e	�h 0����m����i��	� � �   �� ��
�� 0�� .�0 �� �� 0筥 .��� p� �����	�H�@e	�h 0����m����i��	� � à  �� ��L.ڜ������ �����L�ۢ ��
�� 0���� 0�0 �� �� 0� �� �� 0��� p� ���	���@e	�	� ����
�� 0���� 0�0 �� �� 0� �� �� 0��� p� �����	���@e	�	� ����L���Lۭ����L9ݭ���L9ݜ������ �����L}ܢ ��
�� 0���� 0�0 �� �� 0筢 .��� p� ���	���@e	�	� ����
�� 0���� 0�0 �� �� 0筢 .��� p� �����	���@e	�	� ����L����L�ۜ������ �����L1ݢ ���� �� 0���� 0�0 �� �� 0筢 .��� p� ���	���@e	�	� ������ �� 0���� 0�0 �� �� 0筢 .��� p� �����	���@e	�	� ����L����L�ܩ���������� �����L�ݢ �� �� �� 0���� 0�0 �� �� 0筢 .��� p� ���	���@e	�	� ���� �� �� 0���� 0�0 �� �� 0筢 .��� p� �����	���@e	�	� ����L?���L?ݭ� .� .筡�� ��iy��i�� Z� �� ��� ����L�̭���L�̀� ���L�� �� ���� ����L߭�
�� 0�� .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0� �m����i��	� � �   �� ��
�� 0�� .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0� �m����i��	� � à  �� ��LHޭ �������L� ���� �� 0� .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0��m���i��	� � �   �� ���� �� 0� .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0��m���i��	� � à  ���L)ߩ � ��� ����m�����m���� � �{�� ��
������8�������c� � � 筫�� N��������x�
������������x�
������
m��������� �  � 筧�� N�L�� ��
��	�	��L�� ��
�� 0�	 .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0�
�m	���i��	� � �   �� ��
�� 0�	 .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0�
�m	���i��	� � à  ���	L��
 �a�� �Ŝ���8���������������� � �>�� � �ŭ��
���	�LZƭ��LƩ
 �#�� �� �ũ������L�����L� � ����� ���L㭡
�� 0� .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0��m���i��	� � �   �� ��
�� 0� .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0��m���i��	� � à  �� �LL� �������L� ���� �� 0� .�0 �� �� 0筢 .��� p� ���	�H�@e	�h 0��m���i��	� � �   �� ���� �� 0� .�0 �� �� 0筢 .��� p� �����	�H�@e	�h 0��m���i��	� � à  ���L-�m�L/��L#�
 �a�� �ŭ�8���������������� � �>�� � ��LƩ<��P��T��'��R��Y��V��X�:��S��B�� �Z�!�<�"�W�#:�$�\�%�>�&��'�(�[�)�U�*`��� �  `� r �� ���r �� ���`�H�e � ��h`�
&�`�
&
&
&�`�
&
&
&
&�`� �����L `�����	� �
�������� ����
����	������` p� %� � � �  � �� �Li�H�' )��$ �,�' )��% �+h@�-@8���`�8���`� ��� � �� ��� � ��8��	��i�	`P�I�	`i��`��e��`� ��`�� �� � �� �`� �`�L��L��L��L��.��/�	��ف�� ����f�ȩ��� � E� E����LE�� `�ȝE�` H� �.�/�`���	����`�� ��� `���.� 瘤	�'��Ff�e��	e��fjff����`L��	�����L�� 瘠�	��F�e��	e��fjf��몥`F�ejf�����`��	
&	
&	e��e	*��`�� �	�� �L�� � � �� � � `�� � `� � H� 8�� ����� h�� `�� 8�� ��� ��� � � Ȋ� `�Q�R�S�T�Qi��QmR�RmS�SMQ)��SmT�TMR`H��� �	�� ��h�L�� � �H�� h`�H�� �	� ��Ȋ��h�L��
�� � �
���������`� 8I�r �H�I�q �hL�� 8I�q � HȊI�q � �h`� �� � !��	`� ����&	*&��������������`&	*��������`� �� � !��`�c���	� �� �
�����	����������`� � `�� `�  I�� ` �0��<��3��?�%#"$�.�/�5�6�����?�����>�A ������`L  L  L  L  ����joy  ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        <f~fff |ff|ff| <f```f< xlffflx ~``x``~ ~``x``` <f`nff< fff~fff << l8 flxpxlf ``````~ cwkccc fv~~nff <fffff< |ff|``` <ffff< |ff|xlf <f`<f< ~ ffffff< fffff< ccckwc ff<<ff fff< ~0`~    ��   �� 00 ���� 00 ��������� TTTtTTT            fff     ff�f�ff >`<| �� 00 ���� 00 ��    �� 00 ���� 00 ���� 00 ���� 00 ��     0   ~           0` <fnvff< 8~ <f0`~ <ff< f ~`|f< <f`|ff< ~f <ff<ff< <ff>f<           0��������  ~ ~   ے��RR� <f     ��   >>     BBZ~<<<      ��     ��         ��  00000000   ��8   8��   ����������p88p�����������a? <~~~~< �`0��0BBZ~<<<   ����      ���~Z~Z~Z~Z��������~f~f~f~f    ��  ��������%%%%%%2 ~f~f~f~f    BBZ~                                                                                                                                                                                                                                                                                �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ɍ& LR�������l�