
''=@>B"**+@%B&<?.-?./#A, A $ ( ) POWER UP ARROWS   POINTS   FREEZE   WALL     C R O S S  H O R D E FABRIZIO CARUSO C L E A R E D GAME OVER           HYPER  HISCORE LEVEL   FINAL POW RNG SPD joy�������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ����L` ��SL:��� � mS�� ���  ��� s� h��U�V ��S��	� �� ���W�X�T�T��L7��� � mS�� �� ��T ��0 s� h� ���  ���� .� h���	�H�@e	�h ��W�XmT���i��	� � à  ���� � mS�� �� ��T ��0 s� h� ���  ���� .� h����	�H�@e	�h ��W�XmT���i��	� � &à  ���TLU��S ��S��	��L�L�� ��Y�Y�� �L�� -��
 b��Z� �Z �� -��
 � ��� �� �q �� G�8�YH�� �h ���  ��� s� h��\�]� �Z�0 ���  ���^�_�[�[��L�¢ �� �q �� G�8�YH�� �h �� ��[ ��0 s� h� ���  ���� .� h���	�H�@e	�h ��^�_m[���i��	� � à  ��� �� �q �� G�8�YH�� �h �� ��[ ��0 s� h� ���  ���� .� h����	�H�@e	�h ��^�_m[���i��	� � &à  ���[L���YLT�L�� �� � �@��	� �@ N�� L�� ��`�a�`� �a�� �
�`���a��L�� �� � JJJJ���	� �L�� �� )���	� � �L���b�b��`�c�c��L	Ĝd�e�e� ��d��LĢ �b
�� ��d�e ��0 s� h� ��c ���� .� h���	���@e	�	� ���b
�� ��d�e ��0 s� h� ��c ���� .� h����	���@e	�	� ��d�L[��eL[��cLK��bL@é  >) �� >) ��` �� �� � �� ��J ���  �� � �L��Lĩ
 ��  �� �� �vLN������ ��  �� �� �LN� �� m��d��c� c�L���  � �� ��2�3LN� �� m2�2� m3�3 ��L��� �ĩL�� ���� ����" -�� �� �� h���	������ ��׭�L��������v�����5����v��	8���� ����v�� ��v�	�8������  �� ����� �� �� �� �� �� N�� �� ����� �� �� �� �� �� N�� �� ����� �� �� �� �� �� N������w�`������������L�Ƣ ���	 �� �� ��� ��0 s� h���	��e��e	�	�H�@e	�h �����m����i��	� � à  ��� ���	 �� �� ��� ��0 s� h���	��eH�e	�h���	�H�@e	�h �����m����i��	� � &à  ���L���L���v�v ��
 b��������-��&�	�%�#��-�2 �ĩ��i��� �����  Ā�� Lĩ �ĭv��&��)��,��/��0��3��6��9��?��8�9���2���+��-�$�-���w���w�����
������LũL�ĩP �ĩ������L�Ȭ��x�������L�Ȭ�����H����������L�Ȣ ��
�� ��� ��0 s� h���	���e	�	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h���	�H�e	�h���	�H�@e	�h �����m����i��	� � &à  ���L�Ǭ�� ��L����`���������x���*��������� �"��� ����	�u��!�
������'�����u������L�ʜ������ �����L�ɢ ��
�� ����� ��0 s� h� ���� �x G� ���� .� h���	���@e	�	� ����
�� ����� ��0 s� h� ���� �x G� ���� .� h����	���@e	�	� ���L���L�Ȣ �� ������������`� ��
�� ��� ��0 s� h� ��� ���� .� h���	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h� ��� ���� .� h����	�H�@e	�h �����m����i��	� � &à  ���L�ɬ����/��
���i��	����� ��
�����i��	��-��
���i��	����� ��
�����i��	����� �� ��������� ����L�˭�
�� ��� ��0 s� h� ��� ���� .� h���	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h� ��� ���� .� h����	�H�@e	�h �����m����i��	� � &à  ��� �L˭� ������������`� ��
�� ��� ��0 s� h� �� ���� ���� .� h���	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h� �� ���� ���� .� h����	�H�@e	�h �����m����i��	� � &à  ���L�˜���������� �����`�ȍu �̩2 ����`�������������� �̩����L�Ĝ1`� �� ��m����i��	�� � ��������� ����Lέ�J
�� ��� ��0 s� h���	��e��e	�	�H�@e	�h �����m����i��	� � à  ��� ��J
�� ��� ��0 s� h���	��eH�e	�h���	�H�@e	�h �����m����i��	� � &à  ��� �LCͭ� ����m����i��	�� � ������������`� ��J�� �� ��� ��0 s� h���	��e��e	�	�H�@e	�h �����m����i��	� � à  ��� ��J�� �� ��� ��0 s� h���	��eH�e	�h���	�H�@e	�h �����m����i��	� � &à  ����L9� ��� }����x�������������������� ���� �ȱ �L�� �� � }����L�Ҡ���Lќ������ �����LТ �
�� ����� ��0 s� h� ��� ���� .� h���	���@e	�	� ���
�� ����� ��0 s� h� ��� ���� .� h����	���@e	�	� ����Lq���Lqϭf)���	����q��� � ������������L�Ң �
�� ��� ��0 s� h� ��� ���� .� h���	�H�@e	�h �����m����i��	� � à  ��� �
�� ��� ��0 s� h� ��� ���� .� h����	�H�@e	�h �����m����i��	� � &à  ����LBР�)�L�ќ������ �����L�Ң �
�� ����� ��0 s� h� ��� ���� .� h���	���@e	�	� ���
�� ����� ��0 s� h� ��� ���� .� h����	���@e	�	� ����L%���L%Ѡ�� ������������L�Ң �
�� ��� ��0 s� h� ��� ���� .� h���	�H�@e	�h �����m����i��	� � à  ��� �
�� ��� ��0 s� h� ��� ���� .� h����	�H�@e	�h �����m����i��	� � &à  ����L�Ѳ ���J���)e�� Y������� ��� �� ͥ�	����8������� ��� �L�� � U� �� b������ ����5��� �� �� � ������� ���  W��� ���	� ���ĩL��������  Ӎ���͠�� ����� �͠�ޢ �� G�� �͠�ͬ������:���x�m����	�oJi�` [Ӭ�� ��������s`�o��2�o��
 U�)�#�!�o�� U� �� � ��
� U�)i�����m��� [Ӭ�����������r`� �lmm����� PI������` �������LMբ�H����������LGբ ��
�� ��� ��0 s� h� ���  ���� .� h���	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h� ���  ���� .� h����	�H�@e	�h �����m����i��	� � &à  ����Ls���L\�L��������'��*��� �� ������������`� ��
�� ��� ��0 s� h� ����x ���� .� h���	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h� ����x ���� .� h����	�H�@e	�h �����m����i��	� � &à  ����Lrլ���� U��K�`�j��j�o���v����j�j��9�`�6� ��-L׭j���G�`�D� ��#�t����u��@�h�=� ��-�Z����v�	��N�L�K� ��#�>����l��U��R� ��2�$�|� �č���� �� ��i|��i�� ��ZL�`�s��r��s� �Ӏ �� ��L5Ԭ��x��������� �����L�ע ��
�� ����� ��0 s� h� �� ���� ���� .� h���	���@e	�	� ����
�� ����� ��0 s� h� �� ���� ���� .� h����	���@e	�	� ����LF���LFע�����������L�آ ��
�� ��� ��0 s� h� ��� ���� .� h���	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h� ��� ���� .� h����	�H�@e	�h �����m����i��	� � &à  ����L؜�����L�٢�����������L�٢ ��
�� ��� ��0 s� h� ��� ���� .� h���	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h� ��� ���� .� h����	�H�@e	�h �����m����i��	� � &à  ����L�� P���L�؜������ �����L|ڢ ��
�� ����� ��0 s� h� ��� ���� .� h���	���@e	�	� ����
�� ����� ��0 s� h� ��� ���� .� h����	���@e	�	� ����L����L�٩ V� ͬ�����q�m��p�l���h��g���� H֬�� ��`������`�����L�ܬ������� ���/L�ܜ������ �����L�۬�� ��
�� ����� ��0 s� h� ���� ���� .� h���	���@e	�	� ������
�� ����� ��0 s� h� ���� ���� .� h����	���@e	�	� ����L����L�ک�m����	�8�������L�ܬ�� �� ������������L�ܬ�� ��
�� ��� ��0 s� h� ���� ���� .� h���	�H�@e	�h �����m����i��	� � à  ����� ��
�� ��� ��0 s� h� ���� ���� .� h����	�H�@e	�h �����m����i��	� � &à  ����L����L�ڜ�� ����Lެ����Lެ���͠�Lެ��x ���� G� Y�0���x ������ Y�0�� Lޭu������������L ެ�� ���/������� �����L�ݬ�� ��
�� ����� ��0 s� h� ���� ���� .� h���	���@e	�	� ������
�� ����� ��0 s� h� ���� ���� .� h����	���@e	�	� ����LG���LGݢ �` �Ȣ ���L�ܩ `������x�m����	�8�������`���m����	�8��������� �����`� ��
�� ����� ��0 s� h� ���� �x�� ���� .� h���	���@e	�	� ����
�� ����� ��0 s� h� ���� �x�� ���� .� h����	���@e	�	� ����LS���LSޜ�����z�����l �ܪ�f��������
��� ������m������	�8�������� Pբ
�� �� � �Ȁ��������	� � �� 7� ��L�`�g��h� Ӎ�����������������)����x���g���g���h����L=㬠�x��L=��m����	�8��������L���H����������L�� ��
�� ��� ��0 s� h���	���e	�	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h���	�H�e	�h���	�H�@e	�h �����m����i��	� � &à  ����L!��H����������L�� ��
�� ��� ��0 s� h���	���e	�	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h���	�H�e	�h���	�H�@e	�h �����m����i��	� � &à  ����L����L
ଠ��L���H������ʭ���L�⭠
�� ��� ��0 s� h���	���e	�	�H�@e	�h �����m����i��	� � à  ��� ��
�� ��� ��0 s� h���	�H�e	�h���	�H�@e	�h �����m����i��	� � &à  ��� ��L�������� �����L�� ��
�� ����� ��0 s� h���	���e	�	���@e	�	� ����
�� ����� ��0 s� h���	�H�e	�h���	���@e	�	� ����L����L�⩌�m����	�r����m����	�)�������x�m����	�r� �Ȭ��x���1LP�`��J���)e�������w�L���L��/��L��w������� ���)
�� ������ m�����������L��8�������L��.�.���.����.��.����/�w��)��m.�� ���) ����i��	���  ���!��m.�����)����	����.���.�������L�� cĭ-�0��Lͬ���x�fL�Ȝ���`��0������L�� �
�� �� ��0 s� h���	��e��e	�	�H�@e	�h ���m���i��	� � à  ��� �
�� �� ��0 s� h���	��eH�e	�h���	�H�@e	�h ���m���i��	� � &à  ���L���L��
 ��z��L ĩx�m��� � U�)i�  ����� �� �Ȣ
�� �� 7�L�� ]��E� ���4�5�28�4��3�5���3�5�2�4�2�3��k�o�q�p��n =é  Vԩ Vԩ �����  ĩ �� �� ��4�5 N�� ��U��  ĩ ��j��  Ĝ���L�� �
���i��	�� � ��������Ly� ��0 s��
 �� �� ��	 �� ���� .� h���	�H�@e	�h ���m���i��	� � à  ��� ��0 s��
 �� �� ��	 �� ���� .� h����	�H�@e	�h ���m���i��	� � &à  ���L�� �� ��	 �� �� � ��i(��i��� ��L�� I� =�L�����u�v�.�/�0���i�g:�������1�	�-�-�t�c��	����� 
�����w�9�#�8�č<�͍;�@�(�?�̍C�ߍB�G�,�F�ƍJ���I�N�)�M�ǍQ�}�P�U�*�T�̍X���W�	�	��L� �	 ��iY��i�	� ����	 ��iY��i�	�&��� �	 ��iY��i�	���ȩ͑� �	 ��i|��i�	� ����	 ��i|��i�	�$��� �	 ��i|��i�	�x��ȩǑ�	L[� =Ü�������� ��������8�p�l���l���
�f� �� ��f�
�� �l8�
�s�o ���
 ��8�q�m�m ��8�
H�� �h Y��m��8�
�
�f� �� ��f�
��m8�
�r 5Ԝ�������� ����� �� V� � �Ģ�؍�����Lx� ��0 s�� ����	�H�@e	�h ���m���i��	� � à  ��� ��0 s�� �����	�H�@e	�h ���m���i��	� � &à  ���L�� ��  �� ��4�5 N���������L5� ��0 s�� ����	�H�@e	�h ���m���i��	� � à  ��� ��0 s�� �����	�H�@e	�h ���m���i��	� � &à  ���L���`������L�� ��0 s�� ����	�H�@e	�h ���m���i��	� � à  ��� ��0 s�� �����	�H�@e	�h ���m���i��	� � &à  ���LB� c� LĢ�Ѝ�����L�� ��0 s��$ ����	�H�@e	�h ���m���i��	� � à  ��� ��0 s��$ �����	�H�@e	�h ���m���i��	� � &à  ���L�� ��  � �� �o�� N�� �� ����i��	�� � ������ ���Lw� ��0 s��" ����	��e��e	�	�H�@e	�h ���m���i��	� � à  ��� ��0 s��" ����	��eH�e	�h���	�H�@e	�h ���m���i��	� � &à  ��� �L��� ����i��	�� � ��������LL� ��0 s��$ ����	��e��e	�	�H�@e	�h ���m���i��	� � à  ��� ��0 s��$ ����	��eH�e	�h���	�H�@e	�h ���m���i��	� � &à  ���L�� � �� �� �n N� ŭo��� ��
 ����� �� ��
 ����� �� ��
 �� �� �o�� N� Iĩ ��
 ����� �L���i��i�i������- ��  >��)�L����L������)
�����L����� ����L�� ��J �� �� ��� ��0 s� h���	��e��e	�	���@e	�	� ����J �� �� ��� ��0 s� h���	��eH�e	�h���	���@e	�	� ���L
��L
� �L���)�L����%�L������)
�����L��� � � ����L�� ��J G� �� ���  ��0 s� h���	��e��e	�	���@e	�	� ����J G� �� ���  ��0 s� h���	��eH�e	�h���	���@e	�	� ���L��� L�� ̀��) ���� �����/���0������ ͭ0��0 �ک�!�!��L��!��L���H�#�$�"�"��L�� �!
�� ��" ��0 s� h���	���e	�	�H�@e	�h ��#�$m"���i��	� � à  ��� �!
�� ��" ��0 s� h���	�H�e	�h���	�H�@e	�h ��#�$m"���i��	� � &à  ���"L���!L����t��t�
�	 �ĩ-�t�2�3 ��k ���� .� Y��L��n�	��n�k�%� �%���
�� �¢
�� �¢ �%��� ����i��	�� � ���'�(�&� �&��L�� ��0 s��" ����	��e��e	�	�H�@e	�h ��'�(m&���i��	� � à  ���& ��0 s��" ����	��eH�e	�h���	�H�@e	�h ��'�(m&���i��	� � &à  ��� �&L>�� ����i��	�� � ���*�+�)�)��L��) ��0 s��$ ����	��e��e	�	�H�@e	�h ��*�+m)���i��	� � à  ���) ��0 s��$ ����	��eH�e	�h���	�H�@e	�h ��*�+m)���i��	� � &à  ���)L� � �� �� �n N��u���-f�� �߀�u � U� �� b��������@������6���x�
�,�u�'�Y� �č,��� �, ��iY��i�� �� ϩ6� Mϩ=� MϩD� MϩK� MϩR� MϜ-�-��-� �- ��i|��i�� MϢ �- ��iY��i�� M��-�̢
�� ���f�1��l�L��m�L��1�5�o �� Iĩ� �ĭv��v� �� LĢ*�0 �­v�� IĜq�p��n�� ͜� Iĭn�
�o�	�L��n�'�.�.���� ��8�.�� ���.�� I� =é
 �����  � I� =�L�婠� �  `� r �� ���r �� ���`�H�e � ��h`�
&�`�
&
&�`�
&
&
&�`�
&
&
&
&�`� ����`� �`��	l � ��ɢ�L`������	� �
�������� ����
����	������` s� ��� � � �  � �� ��L#�H�' )��$ �0�' )��% �/h@�1@8���`�8���`� ��� � �� ��� � ��8��	��i�	`P�I�	`i��`�L����e��`� ��`�� �� � �� �`� �`�L��L��L��2��3�	���ŀ� ���� �ȩ���� � �� �����L5�� `�ȝ5�` 8� �2�3�`�� ��� `�  ����$L��`���.� ����	�'��Ff�e��	e��fjff����`Lu��	�����L�� �����	��F�e��	e��fjf��몥`F�ejf�����`��	
&	
&	
&	8�H�I�e	�h`��	
&	
&	
&	eH�e	�h`� I�iH�I�i �h`�� �	�� �L��� � � �� � � `�� � `� � H� 8�� ����� h�� `�� 8�� ��� ��� � � Ȋ� `�A�B�C�D�Ai��AmB�BmC�CMA)��CmD�DMB`�H� �h� ȵH� �h� `��  ���� ����  ����	L$�H��� �	�� ��h�L��� � �H�� h`�
�� � �
���������`� 8I�r �H�I�q �hL~�� 8I�q � HȊI�q � �h`� �� �� $���	`� ����&	*&��������������`&	*��������`� �� �� $���`�S���	� ���
�����	����������`� � `�� `�  I�� ` �0��<��3��?����%�&�����/�����.�1 ������`L  L  L  L  ����joy  �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        <f~fff |ff|ff| <f```f< xlffflx ~``x``~ ~``x``` <f`nff< fff~fff << l8 flxpxlf ``````~ cwkccc fv~~nff <fffff< |ff|``` <ffff< |ff|xlf <f`<f< ~ ffffff< fffff< ccckwc ff<<ff fff< ~0`~    ��   Z$f�$$  Z$fY   �� f�$$          $ � $$      $>`<|     Z$f      Z$$f�$$*w* ������� Z$f�$$  Z$fY<~����~<?B��   
	  p �"%�P<fnvff< 8~ <f0`~ <ff< f ~`|f< <f`|ff< ~f <ff<ff< <ff>f< JJJJJJd ***:***    ?@��   $fY    $f   � P� $$       p     P�$$                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ɍ& L���C���&�