����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ����L` Y� 0� ҭ_)� 0���	� �r�:�_)�� 0���	��q�"�_)�� 0���	� �	 0���	��8�� 0� ��L���� 8ĩ�U �ɜh��8��`���a����i�U�_ [Ɯ������ �� ��i���i�� �����Ģ �Щ`� �� C��� "Ŝ���������� Kŭh�
�Ģ PӪ�` Y�  C�LB� =� �� �q �� Y��  W� �� =� Y� 2���	�� �� �� �� Y� �� ��L8¢ ȱ �	q �� r� Y��  W�0 �� =� Y�
�  W��� v� =��	�H�@e	�h Y�� �q �� �q i��	� � Ġ  �� �� �	q �� r� Y��  W�0 �� =� Y�
�  W��� v� =����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q LP� ���r � � 2���	� ���L�L�� Y� F� �� �� �L��� ��
 �� � � � C� ��
 V� � =� �� �q �� -�8�� H�� �h Y��  W� �� =� Y�� � �0 ��  �� Y� �� ��L�â �	� �q �� -�8�� H�� �h r� Y��  W�0 �� =� Y��  W��� v� =��	�H�@e	�h Y�� �q �� �q i��	� � Ġ  �� �	� �q �� -�8�� H�� �h r� Y��  W�0 �� =� Y��  W��� v� =����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q L�� ���q Lb�L�� C� � �@��	� �@ 4� L�� C� � JJJJ���	� �L�� C� )���	� � �L�� F� �� ��Lũ � ��L� F� � �� � �� ��L�Ġ� � 
�� Y� ��0 �� =� Y��  W��� v� =��	���@e	�	� ���� 
�� Y� ��0 �� =� Y��  W��� v� =����	���@e	�	� �� S�L\� ���r LJĠ�q L?�L��  >) �� >) ��` Y� W� 2� � -�J C��  C� 2� �L��  > C� )�!�Ģ �������t���2�^��eL�Ų )� �Ģ �������s���2�^��e�^� )� �Ģ �������v���2�]��e�8� )��Ģ �������u���2�]�e�� ) ��i�	����hL��W���V��#�Z���Y�X��q�r Y�Y�Z ��L/��@`�Y��Z� � ��Y8��Y��Z`�Y�Z` =� � ��� �  ��i���i�� ���r ��L�� =� �� �  ��i���i�	���� � ��r � � � ��֩L�� C� =� � �� �L�� =� � �� Y� �� ��L�Ǣ ȱ �q �� r� Y��  W�0 �� =� Y��  W��� v� =��	�H�@e	�h Y�� �q �� �q i��	� � Ġ  �� �� �q �� r� Y��  W�0 �� =� Y��  W��� v� =����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q L�� ���r L��L�� C� =� � �� �L�� =� �� �� Y� �� ��L�Ƞ� � 
�� Y��  W�0 �� =� Y� �� �q �� Y��� v� =��	�H�@e	�h Y�� �q �� �q i��	� � Ġ  ��� � 
�� Y��  W�0 �� =� Y� �� �q �� Y��� v� =����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q L�� ���r L��L�� Y� F� 2���	�
�� 2���	�
��� � ��L�ɩ � ��� J�	��	�� � 	j� 2� �Р� )�� )�q �� �q �	�r�� )�q �� �q �	�8�� F� � �� � �� �7�� � S�� ���r L&��q L�L�� F�  C�l�	��JJ�U�o��l�p� �� ��d�3�q ���	� 

��� �  ��iE��i�� Y�� ��3 C� C� C񩃢 �Ҡ� �  ��iE��i�� �Р�q ��� �� ��L˩ �� ��L�ȱ ��
�� ��Lˢ �U� �`�^�  ��i���i�� Y�� � 
���� Y� �� Y� S� C�� � 
���� Y� �� Y� S� C� C�w��(�  ��i���i�� Y�8��  C� C�: C�y� ���r � ��q LQ���q LEʩ � �� ��m��� ��\� �  ��i���i�� Y�� �  	� Y� ��) -� C�� �  	� Y� ��) ;� C�  C�x� ���r � ��q ����q ���e� Y�
 C� C� C�z� �ΩТ Y�
 C� C�  C�z� �Ωڢ Y�
 C� C�  C񩄢 �Ωy� Y�
 C� C�  C�~� �Ω�� Y�
 C� C�  C񩈢 �Ω� Y�
 C� C�  C񩉢 �Ω� Y�
 C� C�  C񩊢 �Ωo� Y�
 C� C�l�� C�|� �ΩĢ Y� �� )�
 �� C� �� )�
 �� C� C�s� �Ω� Y�
 C� C�  C񩅢 �Ω� Y�
 C� C�  C񩆢 �έm��%� Y� C�
 C� C񩂢�@�n��l�9�%� Y� C� C�: C񩂢 �ҩ � Y�  C� C� C񩁢 �ҩ� Y�
 C� C�  C�{� �Ω*� Y�  C� C� C�{� �ҩĢ �Щ�� Y�  C� C� C�{� �ҩ`� Y� C� C�l

i C�}� ��L��� W� �� C� ��� �� �	� 8�
i�D�
 W�DJ -�BL��� W� ��� �������� �`�� `���� ��-�� W� ��� ����� W� ��� ���� �`�``�� W� ��� ��L?�� W� ��L����� ��-�� W� ��� ����� W� ��� ���� �`�`` Y� ���  C��  C��  C� 2� �Ҡ 2� fԠ 2� �ժ��L�� Y� 0���	��L�� =� 2���	� � �� Y� �� ��L�Ϡ� � 
�� Y��  W�0 �� =� Y�	�  W��� v� =��	�H�@e	�h Y�� �q �� �q i��	� � Ġ  ��� � 
�� Y��  W�0 �� =� Y�	�  W��� v� =����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q L� �� 0���	� L�� F� � �� � �� ��L�Р� � 
�� Y� ��0 �� =� Y��  W��� v� =��	���@e	�	� ���� 
�� Y� ��0 �� =� Y��  W��� v� =����	���@e	�	� �� S�L�� �� 0���	��L�� Y�?�& 0���	� C� 2���	�� C�Ģ  Ӫ�� ���� L�� Y� =� 2� %���	� � �� Y� �� ��L Ҡ 2���	� �
�� Y��  W�0 �� =� Y� 2���	�� W��� v� =��	�H�@e	�h Y�� �q �� �q i��	� � Ġ  �� 2���	� �
�� Y��  W�0 �� =� Y� 2���	�� W��� v� =����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q L� ��L�� Y� F� � �� � �� ��L�Ҡ 2���	� �
�� Y� ��0 �� =� Y� 2���	�� W��� v� =��	���@e	�	� �� 2���	� �
�� Y� ��0 �� =� Y� 2���	�� W��� v� =����	���@e	�	� �� S�L� ��L�� Y� 2���	�� �� 2���	�� ��� 2���	�� �� 2���	 0��Ȋ�L�� Y� 0���	�� ��� � 0���	��� �� ���� L�� Y� 0���	��. 0���	���! 0���	��� 0���	����� ���� L���LE� Y� 0���	���Z 0���	� C� 2���	�� C񩰢 Y� �ժ�/�mS�S��T 0���	�	8�U� 0���	��� 0� ��L�� C��  C��  C񩈢 Y� �ժ�6��  C��  C񩰢 Y� �ժ��� ����� ������� �� L�� Y� F� 2���	� W� �� Y� � e� ;�8��� � 2���	�� W� �� Y� � e� ;�8�� ��  C��  Ԫ� 2���	�� �� 2���	� ��L�� Y� 0���	� �� x׭���L�� =� � ��L�բ �  ��i���i�� ҭU)�2� �  ��i���i�	�8��� �  ��i���i�	��8��.��  ��i���i�	�r�� �  ��i���i�	��q��r L
� �� 0���	�y��ȩ��U ��L�� C� =� � � � �� �1��  C��  C� ��� �  �� =�  Ӫ�� ��r �ÊL�� Y� 0���	� ��
�7 0���	�� ��B�% 0���	�� W�BmD�� -� j�0�� ���� L�� ���
�'���>�� W�8�>H�� �h j�� �`� �`�` C� =� �� �� Y� �� ��Lrנ� � 
�� Y��  W�0 �� =� Y��  W��� v� =��	�H�@e	�h Y�� �q �� �q i��	� � Ġ  ��� � 
�� Y��  W�0 �� =� Y��  W��� v� =����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q L�� ��L�� C�: C� C�S�TLX� =� �| �� Y� �� ��L<ر  W�0 �� ���	�H�@e	�h Y�� �q �� �q i��	� � Ġ  ���  W�0 �� �����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q L�� �� =� �w �� Y� �� ��L�ر  W�0 �� ���	�H�@e	�h Y�� �q �� �q i��	� � Ġ  ���  W�0 �� �����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q LQ� �� =� �s �� Y� �� ��L�ٱ  W�0 �� ���	�H�@e	�h Y�� �q �� �q i��	� � Ġ  ���  W�0 �� �����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q L�L�� C�  C� C� �iLX© C�  C� C� ��LX©	 C�  C� C� �ULX© C�  C� C� ��LX© C�
 C�ˢ� �� C�
 C� C� ��LX©
 C�â�L"ũ
 C񩇢�L"ũ
 C񩝢�L"ũ
 C񩱢�L"� '۩ C�&�� "ũ  C���� �ک C��� "ũ
 C�E�� "ũ C���L"ũ
 C񩒢�L"� Y� C��  C� C� 2� X�L�� Y�
 C� 2� ��L��
 C�6�� "ũ C���L"� '۩ C񩺢� "ũ
 C�b�� "ũ C�T�� "ũ C�|�� "ũ C񩧢�L"ũ C�p��L"ũȍv�w���l�m��Ѝ����������詼�������������������� ���������	�
��X��`��k���j��u��t�����~����Ǎ�����ʍ�����؍���������������������(������` 8� Q� � 8�L�ڭ=�� *�9�<�� *�8�8��9���7` 2�E� ����� �� � � 8ĭ��� �� � 8ĩ�g�S�T��������U�=�< [΍l ΍o �͍m G΍n i΍p�V�W�h�Y�Z�:��?�<�Y�f�d�@�A � �j�i 3۩2�]�^�`8�q�m���r ƍ��� 8� �� 8ĭ�JJJ�;�l� �� 8� �� �� � 8ĩ  C� C� �Ʃ  C� C� �Ʃ  C� C� �ǩ C�  C� �� �� �� �� x� �� �� �� ��LV� Kŭ?��� C�� C���� Y�X� ��L�� =���	���� � �� Y� �� ��L�ޢ ��
�� Y��  W�0 �� =� Y�� W��� v� =��	�H�@e	�h Y�� �q �� �q i��	� � Ġ  �� ��
�� Y��  W�0 �� =� Y�� W��� v� =����	�H�@e	�h Y�� �q �� �q i��	� � !Ġ  ���q L�� �� 2� 
�S�T Y�g W��� v� j��	�g�� �� ��f�m�@��j��b�	��2�`���2�č1�2 t������0�U��)�1�2 Y�V� ) ��i���i�� Y�V)
 ���Y�(�Z�#������� �� ��i���i�� ������b� �筅���� �������� �� ��i���i�� ������y� �o� �e� �f� Y�d� ��Т �ڢ �� �?� Y�Y� ��<�"�� � ��8���� �7��� �=�O�� �@� Y�Z� ��9�5�� �A� Y�[� ��A��V)��mS�S��T x� 5�Ģ PӪ�P�?�N�� C�� C񩈢 Y� �ժ�0�� C�� C񩰢 Y� �ժ��Ģ �ժ��p�	 P֪� �ӭV)� [ƭV)�p ƍ����
 C� W�DJ -� C�D �ǭp�J� ��JJJJ�� Y�V�W Y��, X� ;�>� C�
 C�> �Ʃ8�> C�
 C�> ���V��W F� � �� ��� �,�� � S�� �����U��l�Lvݭb��l�Lvݭ��W��0�č/����s�� !کdmS�S��T��U�l� -�����<�=J��b��<�:m=�=���^�_�_��@������1� �� ��i���i�	���� �� ��i���i�� ������_����0�`�/�������/�0 �ȭ��
����L�ܭ��� q� � 8� 9� � 8ĭS�T �� ŭS8����T���LM��LMܭT���S��LMܩ'�s�=�t�@�u�>�v�B�w�"�x��y�!�}�,�z�|�$�~�.�{���<�:��:������#���A���'���?���!���B���"��` Y� 2���	�� 0���	����� 2���	� �r��3� 2���	�� 0���	� ���� 2���	� �8������L�� Y� 2� Ҡ �� 2� ��� 2��� Y� 2��� �L�� Y� 2� Ҡ 2��� Y� 2��� ��� �� 2� �L�� C� ��)� ��� �� 2� v�� �� 2� �� 2� ��L�� =��JJJ C��� ��<�\�q ���	� i��	8�� H� � �hi\��i�	�8� ���q ����\�]L�� Y� =� � ��w� �  ��i���i�	����A�A�V)�: ��8�������)�'� ��� �  ��i���i�� Y�� ��\ ��� �  ��i���i�� ���r ��L�� Y� 2���	��& 0���	��� 2���	� � 0���	�8��L�נּ�� �������� ��������� �����` Y� 0���	� �� x�L�� Y� 0���	��� 0� f� 0� �ժ��L��mS�S��T 7Ʃ�f�md�d` �婖�l�m` ��������`��i �٩mS�S��T` ��ȍv�w`� �� ��d ��mS�S�mT�T�N� ����` Y� 0���	����_�� C�� C� 2�  Ӫ� 0� %� �� 0� c�d 0���	� C� 2���	�� C� 2� q� 2�	 �� �΀/ 0� %�� �� � 0� y� 0���� %� -��Ȋ�L�� �� ��L�� ���x����`����<�7L�٩�?�x�Y` ��3������` �� �� ������� `��@�N� �	�
���Z` =��A�=�N� �����[� ��8� �  ��i���i�	�����  ��i���i�	�yȑȩ��r ��L�� F��,��*��+�� �� �� �� ���	��0�`� 0� ��i���i�0��/L��j�G�l��]�0�^�+�U��$�l�%�V�W Y�� Y�ʭ� z� /� j���j`�]�^` e�[�\ ��8�[���\�!��@��V)��Ģ Y�`� Y� ��`� �Ъ�L��`�W���V�@��q�r Y�Y�Z ��L/���`�h�*���%�i� �i �٭e�_������������h������� 5ꩃ�L��` Y� 0� v� 0� B�L�� Y� 0���	���K� 2���	� C� 2���	�� C� 2�  Ӫ�#�
mS�S��T 0� �Ԡ 2���	� ��L�� Y�  C� ��#� ��� �  ��i���i�� ���r � ��L�� Y�j�[�b�V 0���	� C� 2���	�� C�`�  Ӫ�0 0���	� �� 7� 5��b��`� ҩ�mS�S��T x�L�� Y� 0� ҭ_�����0��!�: 0���	� �r�( 0���	��q� 0���	��	 0���	� �8��L�� Y� 0� �� 0� PӪ�L�� 0���	���L�� 0���	� �� 0� ҭm�# 0���	���m 0���	���
�^�'�-�W�n��l�M 0���	��� 0���	�����'��%��# 0���	�� 0���	�����"�� � ��o��l�L�� 0���	����L�� =� � ��r� 2���	��� ��3��T� �  ��iE��i�	���=� �  ��iE��i�	� ���:��  ��iE��i�� ҩmS�S��T x��r �� �� 0���	� C� 2���	�� �ր 0� ��L��,�*�*� ҭ/�0 Y�*� Y� ��*� �Щ*�L��` Y� 0���	� �� 0� ҩ2mS�S��T x��: 5�L��V� )�8�� W�km;�� j���� W�k8�;H�� �h j�� �`�� `�"�S� � ҭ ��� �k�!�&�V)��  ����� ��!� Y�Ţ � � �Щ � �Ъ�L��`�'�W�%� ҭ%����%�k�&�(�V)��% �����%���&� Y�Ţ �%� �Щ%� �Ъ�L��`�m��
�kL��n��l�`��k ���kLT�U���o��l�` =� � ��L/� �  ��iE��i�	���L'� �  ��iE��i�� �Ъ� �� ��)�-� �  ��iE��i�� Ң �  ��iE��i�	��8��� �  ��iE��i�� �Т �  ��iE��i�	����B� �  ��iE��i�� Ң �  ��iE��i�	� 

�� �  ��iE��i�	����r LI�L�褐� �  `� r �� ���r �� ���`� q � HȊq � �h`�H�e � ��h`�
&�`�
&
&�`�
&
&
&�`�
&
&
&
&�`� ����`� �`��	l � ��آ�L`�؅��	� �
�������� ����
����	������` �� �� � � �  � =� ��L	�H�' )��$ ��' )��% �h@�@8���`�8���`� ��� `� 8�� �`�`�  ��	�E�L#�`� ��� � �� ��� � ��8��	��i�	`P�I�	`��e��`� ��`�� �� � �� �`� �`�Le�Le�Le�Le�Le����	������ �����ȩ��� � � ����L5�� `�ȝ5�` 8� �����`���	����`�� ��� `�� �`��� �`��0�� �`�� �`��� �`�ۢ �*`�  ���$L#�`���.� 1�	�'��Ff�e��	e��fjff����`L���	�����L��� 1��	��F�e��	e��fjf��몥`F�ejf�����`��	
&	
&	eH�e	�h`��	
&	e��e	*��`� I�iH�I�i �h`�� �	�� �L�� � � �� � � `�� � `� � H� 8�� ����� h�� `���	����LY�� 8�� ��� ��� � � Ȋ� `�A�B�C�D�Ai��AmB�BmC�CMA)��CmD�DMB`��  #�� ���  #��	Lg�Fj�`H��� �	�� ��h�L�� � �H�� h`�
�� � �
���������`� 8I�r �H�I�q �hLd� 8I�q � HȊI�q � �h`� �� 1� g��	`� ����&	*&��������������`&	*��������`� �� 1� g��`�S���	� ���
�����	����>�����`� � `�� `�  I�� `THE END LURE THE ENEMIES DESTROY MISSILES USE THE JOYSTICK FABRIZIO CARUSO KILL THE SKULL INTO THE MINES MISSILE BASES THE SKULL AND CROSS CHASE FOR POINIS EXTRA LIFE PRESS FIRE GAME OVER AND ITEMS YOU LOST SHOOT AT YOU WON LEVEL    joy �0��<��3��?����%�&�����/�����.�1 ������`L  L  L  L  ����joy  �����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        <f~fff |ff|ff| <f```f< xlffflx ~``x``~ ~``x``` <f`nff< fff~fff << l8 flxpxlf ``````~ cwkccc fv~~nff <fffff< |ff|``` <ffff< |ff|xlf <f`<f< ~ ffffff< fffff< ccckwc ff<<ff fff< ~0`~    ��   �� 00 ���� 00 ��<<<~ZBB�B�����~        <B��Z$$<<B����B< <B��f$>`<| �� 00 ���� 00 ��$f�$f�� 00 ���� 00 ���� 00 ���� 00 �� <f��z$ �~����   8  0<fnvff< 8~ <f0`~ <ff< f ~`|f< <f`|ff< ~f <ff<ff< <ff>f<   ��    �??�     �   <f�$f,�n(($ � $f4v� <Z��Z<�B�����~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ɍ& L����)����