 ,ɲ JJJJ���	� � �L�� ,ɲ )���	� � �L�ǜi�i�� �j�j���i ,ɭj ���j���i��`�  >) �� >) ��` Bɩ @ɠ 1� 1� G�J ,ɠ�  ,ɠ 1� �L�ǩ  >�k)�<����5�� ,ɭ�8� ����#��� 7����� ����������� L���k)�9����2�� ,ɭ� ����"��� 7����� ����������:L���k)�8����18� ,ɭ� ����"��� 7����� ����������� �_�k)�4����- ,ɭ� ���� ��� 7����� �������� ���$�k) �������� ����	��`��`��` ,ɠ�  ,ɠ�  ������  ,ɠ�  ƌ���� L�ǭ������x��m�` Bɭ��� ��LIʢ�p` ,ɭ��L��� )���&��.��8��=��F��P��Z�s� Zɩ ,ɀX� Zɩ ,ɀL� Zɩ ,ɩ�>� Zɩ�0� Zɩ ,ɩ
�(� Zɩ
 ,ɩ�� Zɩ ,ɩ
�� Zɩ
 ,ɩ ,ɩ ,ɩ� Y�L�� B� /ȅ�	� ,ɠ 1ȅ�	�� ,ɩB � /ȅ�	� �� �΃ /� 7� ��L�� B� /� ����������	 Xɭ� �L�� Bɠ � �ɲ ,ɠ� ,ɩ� Bɩ j��l���5�l��.�m������ �l ��i��i�	� ��� ���� ��� �L�ǜm�m���� �m ��i���i�� ��m��` ,ɜn� �n� �K�n ���q ���q �	� ��-��  ,ɠ�  ,ɭn ���q H��q �h ����� �n��n��� L�ǭ����� � ���8����Έ`����`�o�o��1� �o ��i��i�	���� �o ��i�i�� ��o��` ,ɜp�p� ��� mp ,ɠ�  ,ɭ" ��p��L�� ,ɜq�q� ���  ,ɠ� mq ,ɭ# ��q��L�ǩ  ,� ,ɩ l��  ,ɩ ,� l��  ,� ,ɩ ��� ,ɩ  ,ɩ ���r�r��t�u�mr�� Bɭr @ɩ @ɭ�� M� uȠ  ʢ �r ��i���i�� Bɬr�u ,ɩ ,ɩ ,ɩ&� Y�� �r ��i���i�� ��r��������������s�r�r�s�� �r ��i���i�� Bɭr ��r�٭s�r�r�
�(� �r ��i���i�� Bɩ  ,� ,� ,ɪ Y��r�� ���� Bɩ
 ,� ,ɩ  ,ɩ� }���� Bɩ
 ,� ,ɩ ,ɩ� }��� Bɩ
 ,� ,ɩ  ,ɩ� }��� Bɩ
 ,� ,ɩ  ,ɩ'� }���� Bɩ
 ,� ,ɩ  ,ɩ!� }��:� Bɩ
 ,� ,ɩ  ,ɩ+� }��D� Bɩ
 ,� ,ɩ  ,ɩ,� }��N� Bɩ
 ,� ,ɩ  ,ɩ-� }��X� Bɩ
 ,� ,ɩ  ,ɩ"� }���� Bɩ
 ,� ,ɩ  ,ɩ� }���� B� �ɢ )�
 �� ,� �ɢ )�
 �� ,ɩ ,ɩ� }��0� Bɩ
 ,� ,ɩ  ,ɩ(� }��&� Bɩ
 ,� ,ɩ  ,ɩ)� }�����g� Bɩ ,ɩ
 ,ɩ ,ɩ%��;���9�g� Bɩ ,ɩ ,�: ,ɩ%� Y��b� Bɩ  ,ɩ ,ɩ ,ɩ$� Y���� ��r�r��+� �r ��iĨ�i�� Bɩ  ,� ,� ,ɩ� Y��r�έ���� Bɩ ,ɩ ,ɩ� ,ɩ���� Bɩ ,ɩ ,ɩ< ,ɩ � Y��� Bɩ ,� ,ɢ �� �Ơ< �� ,ɩ � Y��� Bɩ ,ɩ ,ɢ �� �Ơ< �� ,ɩ � Y��� Bɩ ,� ,ɢ �� �Ơ< �� ,ɩ �LY��)�t����	8�t���
�� @ɭ�J Gʍ�`�)�u����	8�u���
 @ɭ�J Gʍ��
��`�)���)���)��� �`�� `������ �`�� `��� *� `�� )���)��	�)��`�`��)�� �`� ` Bɠ Zɠ�  ,ɠ�  ,ɠ�  ,ɠ 1� Y�� 1� �L�ǜv�v��1� �v ��i�i�� Bɭv ,ɩ ,ɩ  ,ɩ� Y��v��`����#���� ���
����������` B� /ȅ�	��'��  ,ɠ�  ,ɠ 1ȅ�	� � /ȅ�	� ���  ,ɠ�  �� /ȅ�	��L�� ,ɜw� �w� �K�w ���q ���q �	� ��-��  ,ɠ�  ,ɭw ���q H��q �h ����� �w��w��� L�� Bɭ��& /ȅ�	� ,ɠ 1ȅ�	�� ,ɩ�� ����� ���� L�� Bɠ � �ɲ ,ɠ� ,ɠ������	� �� ��� �L�� B� /ȅ�	� ,ɠ 1ȅ�	�� ��L�� Bɠ� �ɠ� ��� ��ȱ � /Ƞ�Ȋ�ȱ �ȱ �L�� B� /ȅ�	� ��� � /ȅ�	���� �� ���� L�� Bɠ � �ɲ������	��� ���� H� ��� �hL�ǜ�L� ,ɠ� �� ��� ��� ���
� �����L�� Bɠ � �ɢ � ;� B� �� Bɢ � d� aƍx�� � ;� B� �� Bɢ � d� aƍy�x ,ɭy ����x��y��� ��� �L�� ,ɠ� � ͇�!� ͆� @ɭ�m��� 4� b�0�� ���� L�� ,ɢ � ���#�� ��� @ɭ�m��� 4� b�0�� ���� L�� Bɠ � �ɭ��O� @ɭ� 4� b�0?� @ɭ��� b��+�� @ɭ� 4� b�0�� @ɭ�m��� b�0�� ���� H� ��� �hL�� Bɠ � �ɭ��O�� @ɭ� 4� b�0=�� @ɭ��� b��'� @ɭ� 4� b�0� @ɭ�m��� b�0�� ���� H� ��� �hL�� ,ɠ�  ,ɠ�  ,ɭ. �L�ǩ  ,� ,ɩ ,ɭ���LN��
 ,ɩ  ,ɭ �� ,ɩ  ,ɭ �� ,ɩ  ,ɭ �� ,ɩ  ,ɭL�� ,ɩ  ,ɩ ,ɢ ��LN�� ,ɩ  ,� ,ɢ �� 4�LN� � �� [� r�L��� ,ɩ  ,ɩ ,ɢ ��LN�� ,ɩ  ,� ,ɢ �LN�� ,ɩ
 ,ɩ��� �� ,ɩ
 ,ɩ ,ɢ �LN�� ,ɩ���Ll��
 ,ɩY��Ll��
 ,ɩd��Ll�� ,ɩn��Ll� ��� ,ɩ$�� l��  ,ɭ� ��� ,ɩ⢱Ll� 0��
 ,ɩ��� l�L[��
 ,ɩN��Ll��
 ,ɩ4�� l�� ,ɩ�� l�� ,ɩ�Ll� Bɩ ,ɠ�  ,ɩ ,ɠ 1� N�L�� Bɩ
 ,ɠ 1� ��L�� Bɜz�{�z8� ��{�� ��H� ,ɩ
 ,ɩ ,ɭz�{ N��m������z�{ �� �� .� ��mz�z���{��L�� ��� ,ɩ ,ɩ�� ��  ,ɩ	 ,ɩ��� �� ,ɩ ,ɩ��� �� ,ɩ ,ɩ� �� ,ɩ ,ɩ! �� ,ɩ	 ,ɩB ��	 ,ɩ ,ɩ$ �� ,� ,ɩ# �� ,ɩ ,ɩ? �� ,ɩ ,ɩ ��
 ,ɩ ,ɩ;L� ��~� ,ɩ ,ɩw�� �� ,ɩ ,ɩ��� ����� ,ɩ
 ,ɩ����� ,ɩ
 ,ɩ��� �� ,ɩ ,ɩ��� �� ,� ,ɩ��� �� ,ɩ ,ɩ ,ɢ � N��	 ,ɩ ,�: ,ɭ� N��	 ,�: ,ɩ ,ɭ��� N�����	 ,� ,ɩ ,ɢ � N��|�	 ,ɩ ,ɩ ,ɢ �| N��}�}�|�
� .��}���|�|�~���ǩ
 .ƭ�� ,ɩ ,ɩϢ�L�`� ,ɩB��Ll����� ������� �����`������ � ���`�����������n������@�#�$������Ѝ������-�.������� K������������	 K��������#�$�
 K������������ K������A�B��x�7�8�� �K�L�x�U�V�}�_�`����������-�.���K���� �ƍ����#�$ �ƍ#�$�� �ƍ��A�B �ƍA�B�K�L �ƍK�L`�����������!������=�����������6�����"�6�!���6�D�5���,�i�+���@���?���J���I���T���S���^���]` 0� �����O� ,ɭ
i ,ɢ �
���i��	��� �� ,ɭ
i ,ɢ � ��i¨�i��� ���� [� 0�L%��������}������� ���|���� *�{�{��|���z` ���E� �ǜ� � � [� 0�������������
������������������ +� l��� -��� A��� 	��� L��� 鉭�%��������	����������	��
�����:��� ����� �� �ƍ����~������,������������ I� ���� R� 끍� 0� ǎ 0��JJ����� f��� 0� �� ވ Z� [� 0��� Ƅ������ K������� h� � C�������� K������ ��L3� ������� ,ɭ� ,ɭ.��� ,ɭ� ,ɭ �	���� � � ��������� Bɭ� @ɢ�� u� bǐ�	�� �� (� T������� ���@��;���
�1� � ��i���i�	���� � ��i���i�� ���� � C� ����� ������ .ƭ���� ,ɭ� ��� .Ʃ� y���� y���� y���� y��� y���� Bɩ�� ��� y��&� y���� Bɩ�� � ��X� y���� Bɩ�� ��{��:� y��z��0� y��}�!�D� y���� Bɩ�� ��|��N� y��� ,ɭ� ,ɩ�� Bɭ� �������*�����"�m������ �� ��i���i�� ���������� 񋭄)��J 끍�����
 ,� @ɭ�J G� ,ɭ� �������
 @ɭ�J G� ,ɩ
 ,ɭ� l� 0�������������L������L���Ln������ ,ɭ� ,ɭ.��� ,ɭ� ,ɭ �	���� � � 0�� @ɩ �� Bɭ� @ɩ �� c� �����4����-�������!��������������	��� 0������ >Ȫ� 0� ��������J������~m������������ K��c���I��	������ �
��
 �Ǎ��% 0�����������������������
���Lܔ��8������������� [� 0� Ӑ [���� H� 0� � [�L���'��=��@��>��B��"����!� �,��.�:��$�!�.��#�<�":�$:�%��&�#�'�A�+�'�(�?�)�!�,�B�-�"�.` Bɠ� �ɠ � �ɠ ��������	��� �r�� ��� �����	���8������H� � ����hL�� B� /� 7� Xɩ�� _��� /��� Bɩ�� _�L�� B� /� 7� /��� Bɩ�� _���
 Xɩ�� _�L�� ,ɠ� �ɥ� @��� ��)� �s�q�� �o�� ͝��	�� �\���
�0�� 7�������	���q��8��	���8���'��
��� 7���	���r���� 욠� �ȱ �L�� ,ɠ� �ɥ� 瞪� ��)� ��s�� 욀q�� p���	�� 욀^���
�/�� 7������	���r��9��	���8���(���
��� 7���	����q��	�� �� �ȱ �L�� ,� ��)� ��
� 1� �� 1� �L�ǭJJJ�0�/�/��;���m/���	�0i��8�/H� � �hi���i�	�8�0��/����/�/����/����/��`���m�1�1���`� �1 ��i���i�	���D ��8������� �1 ��i���i�� Bɬ1�� �� �1 ��i���i�� ��1���1�1���a� �1 ��i���i�	���D ��8������� �1 ��i���i�� Bɬ1�� ��� �1 ��i���i�� ��1��` B� /ȅ�	�� @ɭ� 4� b�0& /ȅ�	�� @ɩ8�H�� �h b��� ���� L�� B� /ȅ�	��
 W�L�� B� /ȅ�	��� *� L�� Bɩ�� ���	 /� ������ *��� /� *���� �L�� B� /ȅ�	� @ɭ� 4� b�0( /ȅ�	� @ɩ8��H�� �h�� b��� ���� L�� B� /ȅ�	���
 W�L�� B� /ȅ�	���� *� L�� Bɩ�� ����	 /� ������� Ϟ�� /� Ϟ��� �L�� Bɠ 1ȅ�	��& /ȅ�	��� 1ȅ�	� � /ȅ�	�8��L�ǭ��� ��I�8m����I�m����-�. ��I�8m-�-�I�m.�.�#�$ ��I�8m#�#�I�m$�$���� �� ��I�8m����I�m���` B� /� 7���� � /ȅ�	� �� �L�� B� /� � /� ����� /� u����L�� �����m������m���`� ���m������n����`�2�2��`� �2 ��i�i�� ����2� �2 �ȅ�i�	�� ,ɢ �2 ��i��i�	�� 덀�2 ��i�i�� 7��2�� ���������`���	��������������	8�i���m�����Lr� ����|����`�3�3�2� ��3��
m���������m��������`��!� � �Ƞ
 ��m����m����N� ��m������ ������ LK� Bɠ � �ɠ��O�� ,ɭ� ,ɥ� ��������� �ƥ� ���v� ,ɠ� ,ɠ���� Bɥ��	 �� ��Q������ �5� �1���� 㟲 ,ɠ� ,ɠ���� Bɥ��	 �� ��ȱ��� 4ǑȊ�� ��� �L�� ���@�#�$`�����z ���LK�������X��X��` W����3�����d�-�.�LK� � �� W���A�B�LK����Ls��5�5��Ls��4�4��Lm�� �4 ��i��i�	���Lg�� �4 ��i⨊i��� $���u� �q� �4 �ȅ�i�	�� ,ɢ �4 ��i��i�	�� ,ɭ  �� .Ƣ �4 ��i��i�	� ��ȩ�� �4 ��i⨊i�� �� .��4L���5L������N� �K�L�d���LK������������ �U�V� K��6�6���?� �6 ��i���i�	���"� �6 ��i���i�� ���m������6��`����������x���}�_�``�~��������_�`� K��������`����_�`�LK� ,ɲ �� �@� ,ɩ  ,ɭ) �� ,ɩ��� l�� ,ɩ  ,ɭ �� ,ɩ� l�� ��� L�� ,ɩc8��7� �� m����
�c����� [�L�� ,ɠ 1ȅ�	���:���! ��8������� Zɠ�  b�� 1� �� 1� Ɋ�� �L�ǭ��V������+���&�� @ɭJJ �� b�0����&���(��� ��������������LK�`΋Ό`�����)�3 ,������8�8�� � �8 ��i⨊i�� Bɭ8
 Ĥ�8�٭�������)?�
������`�8��8�8���� �8 ��i���i�	���ݭ8���2�� �8 ��i���i�� Bɭ� ,ɭ� ,ɩ ,ɩ� Y�L��`�������а�m�` Bɭ��� ��LIʢ�@` ,�����������` Bɠ � �ɲ ,ɠ� ,ɩ� Bɩ j��9���Y�9��R�m������ �9 ��i��i�	� ���9 ��i�i�� 7������	�� U���8��� ��� �L�ǜ:�:��� �: ��i⨊i�� d��:��`�;�;��1� �; ��i��i�	���� �; ��i⨊i�� ��;��` Bɠ � �ɲ ,ɠ� 덩 ����������2m����� ��� 7�� ��� �L�ǜ<� �<�� ��ią�i�	�����<`� �<�ک` ,ɢ �  ��ią�i�	���<� �  ��iĨ�i�� Bɠ� ��� F�� �  ��iĨ�i�� Bɠ� ��� �L�ǭ�)��=�=�� E��=��=�=�� ϧ�=��`�������`�������������8�����>������8�������������?�> ,ɭ? ୪�]� �� ��i��i�	�>�� �� ��i��i�	�?��� �� ��i��i�	�ȑ� �� ��i�i�� �����` ,ɠ 1ȅ�	������ 1� ��� Zɠ�  ��L�ǜ@�@��"� �@ ��iĨ�i�� Bɬ@�� ��@��` Bɠ � �ɠ��L��� 1ȅ�	� ,ɠ 1ȅ�	�� ,ɥ� ����L��� 1� 7�� 1ȅ�	� ��������� ���m����L���L����	���8����� ��A��J�A�L���L���� 7��� Bɠ�  ���� ����� ,ɠ� ����� ,ɠ� ƌ��C�m������� ��� ,ɠ� 덭��������� Bɭ� � � ����� ��AL�� ��� �L�� ,ɜB�B���=� �B ��i���i�	��� � Zɠ�  ,ɢ �B ��i���i�� p��B��L�� Bɠ� �ɠ � �ɠ��y� ,ɠ� ,ɥ� ����c� ,ɠ� ,ɠ������	� �� ���� 7�� ��� � P�������	�� U����	���8����� �� � � ����L�� BɜC�C��4� �C ��i��i�	��� Xɢ �C ��i⨊i�� ���C��L�� ,ɠ� �ɥ� 7�� � �
���� �)��	���r�'��	��Șq���	��Ȁ��	���8���� �ȱ �L�� ,ɠ� �ɠ��Lg��� ����!� ,ɠ� ����� ,ɠ� ƌ��Lg�� ��������G���
�B�i�=�g��2���0��������i��g���������d�	�b� ߯����o�D�D��d��D�u�U� �D ��i���i�	���=� �D ��i���i�	� ��~��D ��i���i�� 7��m����� ��D��� ,ɠ� � � ����� Bɠ�  ߫�� ��� �ȱ �L�� ,ɲ ����#��0� 1ȅ�	��8��.� 1ȅ�	��� 1ȅ�	� �8��� 1ȅ�	� �q�L�� ,ɜE� �E��Q �ȅ�i�	�� ��� �5�E ��i��i�	� �� ��E ��i��i�	ȱ���� ���E���L�� ,ɭ��Lܯ� �  ��ią�i�	���Lܯ���Lܯ����Lܯθ [�� ������ �  ��ią�i�	�������1� �  ��ią�i�	��8�����\�� ,ɭ� ,ɩ@ ��I���.��  ��ią�i�	������)�� ,ɭ� ,ɩ> ��� �  ��ią�i�	�������3� �  ��ią�i�	��8������c�� ,ɭ� ,ɩ' ��P����1� �  ��ią�i�	�������+�� ,ɭ� ,ɩ= ��� �  ��ią�i�	����� �  ��iĨ�i�� ���� �  ��iĨ�i�� Bɭ� �L�� B� /ȅ�	� �� /� 7��m����� ��~ P�L�� ,ɢ �  �ƍG�H�F�F��L���� � 
�� BɭF @ɩ0 �� c� Bɠ�  @ɢ�� u� cƅ�	�H�@e	�h BɭG�HmF���i��	� �  ��  ʠ� � 
�� BɭF @ɩ0 �� c� Bɠ�  @ɢ�� u� c����	�H�@e	�h BɭG�HmF���i��	� � ��  ��FL"�L�� ,ɜI�J�J� ��I��L���� � 
�� BɭI�J Bɩ0 �� c� Bɠ�  @ɢ�� u� cƅ�	���@e	�	� ���� 
�� BɭI�J Bɩ0 �� c� Bɠ�  @ɢ�� u� c����	���@e	�	� ��I�L��JL�L�ǩ�� �  `BEFORE   TO UNLOCK SECRET LEVEL FOUND USE THE JOYSTICK DESTROY MISSILES KILL THE SKULLS KILL ALL SKULLS FABRIZIO CARUSO KILL THE BOSS CROSS SHOOT PRESS FIRE EXTRA LIFE GAME OVER YOU LOST HISCORE  YOU WON SECRETS VICTORY THE END SCORE ITEMS LEVEL OF  B !  . - " ENEMY   SKULL   BOSS    BULLETS POWER   MINE                 SECRET FOUND joy������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ����L` BɜSL:��� � mS�� Bɠ�  @ɩ� �� cƍU�V /ȬS��	� �� �ƍW�X�T�T��L7��� � mS�� �� BɭT @ɩ0 �� c� Bɠ�  @ɢ�� u� cƅ�	�H�@e	�h BɭW�XmT���i��	� �  ��  ʠ� � mS�� �� BɭT @ɩ0 �� c� Bɠ�  @ɢ�� u� c����	�H�@e	�h BɭW�XmT���i��	� � ��  ��TLU��S /ȬS��	��L�L�� BɜY�Y�� �L�� Xɩ
 �ʍZ� �Z [� Xɩ
 p� &ʢ �� �q �� 4�8�YH�� �h Bɠ�  @ɩ� �� cƍ\�]� �Z�0 �Ǣ  �ƍ^�_�[�[��L�¢ �� �q �� 4�8�YH�� �h �� Bɭ[ @ɩ0 �� c� Bɠ�  @ɢ�� u� cƅ�	�H�@e	�h Bɭ^�_m[���i��	� �  ��  ʢ �� �q �� 4�8�YH�� �h �� Bɭ[ @ɩ0 �� c� Bɠ�  @ɢ�� u� c����	�H�@e	�h Bɭ^�_m[���i��	� � ��  ��[L���YLT�L�� ,ɢ � �@��	� �@ BǢ L�� ,ɠ�  @ɠ�  @ɩ� �� cƍa�b�  �� �ƍc�d�`�`��L�à� � 
�� Bɭ` @ɩ0 �� c� Bɠ�  @ɢ�� u� cƅ�	�H�@e	�h Bɭc�dm`���i��	� �  ��  ʠ� � 
�� Bɭ` @ɩ0 �� c� Bɠ�  @ɢ�� u� c����	�H�@e	�h Bɭc�dm`���i��	� � ��  ��`L�L�ǭ�� )�8�� @ɭ�m��� b���� @ɭ�8�H�� �h b�� �`�� `�d�S�b� 7��b���b���c�&��)��b �ê����b��c� Bɩ�� _��b� ��b� Ɋ��L�`�i�W�g� 7��g����g���h�(��)��g �ê����g���h� Bɩ�� _��g� ��g� Ɋ��L�`����
��L�ĭ�����`��� �ĩ��L4ĭ������`�e�e��`� �e ��i���i�	���L(Ƣ �e ��i���i�� Ɋ�� � �ɢ )�/�e ��i���i�� 7�� �e ��i���i�	��8��� �e ��i���i�� �� �e ��i���i�	����d� �e ��i���i�� 7�� �e ��i���i�� Bɢ �e�� Bɩ @ɭ�� M� uȠ  ʢ �e ��i���i�	����eL"� ,ɜf�f� �#�g�h�h���g��
�g���h���f��L�Ǣ r �� ���r �� ���`�H�e � ��h`�
&�`�
&
&�`�
&
&
&�`�
&
&
&
&�`��	l � ����L`���˅	� �
�������� ����
����	������` �� �Ʃ � � �  � �� ��L�H�' )��$ �L�' )��% �Kh@�M@8���`8���`�8���`�  �ɦ	�E�Lɥ`� ��� � �� ��� � ��8��	��i�	`P�I�	`i��`��e��`� ��`�� �� � �� �`� �`�LzƠLzƠLzƠLzƠLzƍN��O�	����� �����ȩǑ�� � � ����L5�� `�ȝ5�` 8� �N�O�`���	����`�� ��� `�� �`��� �`��0�� �`�� �`��� �`�ۢ �*`�  �ɥ�$L�`���.� ɘ�	�'��Ff�e��	e��fjff����`L�Ȇ	�����L�ȅ ɘ��	��F�e��	e��fjf��몥`F�ejf�����`��	
&	
&	eH�e	�h`� I�iH�I�i �h`�� �	�� �L�Ǡ � � �� � � `�� � `� � H� 8�� ����� h�� `�� 8�� ��� ��� � � Ȋ� `�A�B�C�D�Ai��AmB�BmC�CMA)��CmD�DMB`�H� �h� ȵH� �h� `��  Ʌ� �ǆ�  Ʌ�	L�ʆFj�`�FjFj�`�FjFjFj�`�FjFjFjFj�`H��� �	�� ��h�L�Ǡ � �H�� h`�
�� � �
���������`� 8I�r �H�I�q �hLyƠ 8I�q � HȊI�q � �h`� �� � �ʥ�	`� ����&	*&��������������`&	*��������`� �� � �ʥ�`�S���	� ���
�����	����������`� � `�� `�  I�� ` �0��<��3��?����%�&�����/�����.�1 ������`L  L  L  L  ����joy  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������        8l����� ������� <f���f< ������� ������� ������� >`���f> ������� �00000� �| ������� ������� ������� ������� |�����| ������� |�����z ������� x��|�| �000000 ������| ����l8 ������� ��|8|�� ���x000 �8p��    ��   �� 00 ���� 00 ��<<<~ZBB�~��~<~�        <B��Z$$<<B����B< <B��f$>`<| �� 00 ���� 00 ��$f�$f�� 00 ���� 00 ���� 00 ���� 00 �� <f��z$�B4,B�  8  Z~Z~Z~Z~<fnvff< 8~ <f0`~ <ff< f ~`|f< <f`|ff< ~f <ff<ff< <ff>f<   ��    �??�   ������ <f�$f,�n(($ � $f4v� <Z��Z<<~��~<~�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        �������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ɍ& L����0����